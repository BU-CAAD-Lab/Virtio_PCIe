parameter PARAMETER_PCIE_CONTROLLER_INST_NUM_QUEUES = 2;
parameter PARAMETER_PCIE_CONTROLLER_INST_SLEEP_TIMER_VAL = 100;
parameter PARAMETER_DEBUG_ADDR_WIDTH = 32;
parameter PARAMETER_DEBUG_DATA_WIDTH = 32;
parameter PARAMETER_DEBUG_CLKS_PER_BIT = 125;
parameter PARAMETER_BRAM_INTF0_ACCESS_CTRL_NUM_PORTS = 4;
parameter PARAMETER_BRAM_INTF0_ACCESS_CTRL_PORT_IDX_BITS = 2;
parameter PARAMETER_ENDPOINT_SELECT_INST_AXI_BUS_WIDTH = 128;
parameter PARAMETER_ENDPOINT_SELECT_INST_AXI_ADDR_WIDTH = 64;
parameter PARAMETER_DW_CONVERTER_DATA_A_WIDTH = 128;
parameter PARAMETER_DW_CONVERTER_DATA_B_WIDTH = 32;
parameter PARAMETER_DW_CONVERTER_ADDR_WIDTH = 32;
parameter PARAMETER_MAIN_MEMORY_ADDR_WIDTH = 14;
parameter PARAMETER_MAIN_MEMORY_DATA_WIDTH = 32;
parameter PARAMETER_MAIN_MEMORY_INITIALIZE = 1;
parameter PARAMETER_MAIN_MEMORY_INIT_FILE = "./cpu_firmware.hex";
parameter PARAMETER_INTF_SPLITTER2_DATA_WIDTH = 32;
parameter PARAMETER_INTF_SPLITTER2_ADDR_WIDTH = 32;
parameter PARAMETER_INTF_SPLITTER2_STRB_WIDTH = 4;
parameter PARAMETER_INTF_CONCAT2_DATA_WIDTH = 32;
parameter PARAMETER_INTF_CONCAT2_ADDR_WIDTH = 32;
parameter PARAMETER_INTF_CONCAT2_STRB_WIDTH = 4;
parameter PARAMETER_CPU_ENABLE_COUNTERS = 1;
parameter PARAMETER_CPU_ENABLE_COUNTERS64 = 1;
parameter PARAMETER_CPU_ENABLE_REGS_16_31 = 1;
parameter PARAMETER_CPU_ENABLE_REGS_DUALPORT = 1;
parameter PARAMETER_CPU_TWO_STAGE_SHIFT = 1;
parameter PARAMETER_CPU_BARREL_SHIFTER = 0;
parameter PARAMETER_CPU_TWO_CYCLE_COMPARE = 0;
parameter PARAMETER_CPU_TWO_CYCLE_ALU = 0;
parameter PARAMETER_CPU_COMPRESSED_ISA = 0;
parameter PARAMETER_CPU_CATCH_MISALIGN = 1;
parameter PARAMETER_CPU_CATCH_ILLINSN = 1;
parameter PARAMETER_CPU_ENABLE_PCPI = 0;
parameter PARAMETER_CPU_ENABLE_MUL = 0;
parameter PARAMETER_CPU_ENABLE_FAST_MUL = 0;
parameter PARAMETER_CPU_ENABLE_DIV = 0;
parameter PARAMETER_CPU_ENABLE_IRQ_QREGS = 1;
parameter PARAMETER_CPU_ENABLE_IRQ_TIMER = 1;
parameter PARAMETER_CPU_ENABLE_TRACE = 0;
parameter PARAMETER_CPU_REGS_INIT_ZERO = 0;
parameter PARAMETER_CPU_MASKED_IRQ = 0;
parameter PARAMETER_CPU_ADDR_WIDTH = 32;
parameter PARAMETER_CPU_DATA_WIDTH = 32;
parameter PARAMETER_CPU_STACKADDR = 16384;
parameter PARAMETER_CPU_LATCHED_IRQ = 16384;
parameter PARAMETER_CPU_PROGADDR_RESET = 0;
parameter PARAMETER_CPU_PROGADDR_IRQ = 16;
parameter PARAMETER_CPU_ENABLE_IRQ = 0;
